magic
tech sky130A
magscale 1 2
timestamp 1730636500
<< locali >>
rect 6660 45044 6774 45076
rect 6660 44996 6692 45044
rect 6740 44996 6774 45044
rect 6660 44962 6774 44996
rect 6686 44176 6746 44962
<< viali >>
rect 6692 44996 6740 45044
<< metal1 >>
rect 14928 45082 15070 45118
rect 6660 45050 6774 45076
rect 6660 44990 6686 45050
rect 6746 44990 6774 45050
rect 6660 44962 6774 44990
rect 14928 45030 14970 45082
rect 15022 45030 15070 45082
rect 14928 44988 15070 45030
rect 15490 45060 15606 45094
rect 15490 45008 15520 45060
rect 15572 45008 15606 45060
rect 2466 44748 2494 44782
rect 14982 44748 15010 44988
rect 15490 44972 15606 45008
rect 16038 45068 16146 45100
rect 16038 45016 16066 45068
rect 16118 45016 16146 45068
rect 16038 44976 16146 45016
rect 17704 45088 17808 45124
rect 17704 45036 17726 45088
rect 17778 45036 17808 45088
rect 17704 45012 17808 45036
rect 18244 45098 18370 45124
rect 18244 45022 18258 45098
rect 18344 45022 18370 45098
rect 2466 44720 15010 44748
rect 2466 25694 2494 44720
rect 15523 44674 15568 44972
rect 2766 44649 2818 44652
rect 3365 44649 15568 44674
rect 2766 44629 15568 44649
rect 2766 44614 3410 44629
rect 2766 29010 2818 44614
rect 16076 44579 16107 44976
rect 2887 44548 16107 44579
rect 2887 29844 2918 44548
rect 17738 44517 17779 45012
rect 18244 44988 18370 45022
rect 18796 45064 18910 45088
rect 18796 45012 18834 45064
rect 18886 45012 18910 45064
rect 3007 44476 17779 44517
rect 3007 40774 3038 44476
rect 18288 44448 18316 44988
rect 18796 44982 18910 45012
rect 27596 45066 27686 45084
rect 27596 45014 27616 45066
rect 27668 45014 27686 45066
rect 27596 44994 27686 45014
rect 3080 44420 18316 44448
rect 18845 44450 18875 44982
rect 25160 44866 25256 44880
rect 25160 44806 25176 44866
rect 25236 44856 25256 44866
rect 27310 44863 27430 44882
rect 27310 44856 27336 44863
rect 25236 44817 27336 44856
rect 25236 44806 25256 44817
rect 25160 44796 25256 44806
rect 27310 44811 27336 44817
rect 27388 44811 27430 44863
rect 27310 44786 27430 44811
rect 19192 44450 19258 44454
rect 18845 44448 19258 44450
rect 18845 44420 19198 44448
rect 2998 35544 3046 40774
rect 2588 28979 2824 29010
rect 2587 28946 2824 28979
rect 2587 28214 2654 28946
rect 2700 28881 2840 28884
rect 2870 28881 2934 29844
rect 2700 28878 2934 28881
rect 2700 28758 2706 28878
rect 2826 28786 2934 28878
rect 2826 28758 2893 28786
rect 2700 28755 2893 28758
rect 2700 28750 2840 28755
rect 2587 28198 2844 28214
rect 2587 28105 2712 28198
rect 2630 28078 2712 28105
rect 2832 28078 2844 28198
rect 2630 28070 2844 28078
rect 2466 25666 2958 25694
rect 2930 24522 2958 25666
rect 2994 24864 3050 35544
rect 3080 25602 3108 44420
rect 19192 44396 19198 44420
rect 19252 44396 19258 44448
rect 19192 44390 19258 44396
rect 27628 44358 27656 44994
rect 3368 44330 27656 44358
rect 3368 32606 3396 44330
rect 30072 34878 30078 34998
rect 30198 34962 30204 34998
rect 30198 34915 30409 34962
rect 30198 34878 30204 34915
rect 3318 32578 3396 32606
rect 3080 25574 3348 25602
rect 3176 24864 3232 24870
rect 2994 24808 3232 24864
rect 3096 24796 3232 24808
rect 3096 24780 3236 24796
rect 3096 24704 3132 24780
rect 3214 24704 3236 24780
rect 3096 24676 3236 24704
rect 2930 24494 3072 24522
rect 3044 22610 3072 24494
rect 3044 22582 3330 22610
rect 29518 20844 29524 20856
rect 29462 20816 29524 20844
rect 5590 18590 5642 18596
rect 2732 18538 2738 18590
rect 2790 18578 2796 18590
rect 2790 18550 5590 18578
rect 2790 18538 2796 18550
rect 5590 18532 5642 18538
rect 2582 18462 2666 18478
rect 2582 18410 2598 18462
rect 2650 18450 2666 18462
rect 4294 18462 4362 18470
rect 4294 18450 4302 18462
rect 2650 18422 4302 18450
rect 2650 18410 2666 18422
rect 2582 18394 2666 18410
rect 4294 18410 4302 18422
rect 4354 18410 4362 18462
rect 4294 18404 4362 18410
rect 29462 17892 29490 20816
rect 29518 20804 29524 20816
rect 29576 20804 29582 20856
rect 27224 17864 29490 17892
rect 27224 17850 27288 17864
rect 27084 17838 27288 17850
rect 27084 17822 27252 17838
rect 29508 17121 29514 17132
rect 29489 17080 29514 17121
rect 29566 17080 29572 17132
rect 11376 16722 11450 16732
rect 11376 16716 11384 16722
rect 10633 16673 11384 16716
rect 7514 16526 7520 16582
rect 7576 16526 7582 16582
rect 7520 16278 7576 16526
rect 7520 16216 7576 16222
rect 10633 15528 10676 16673
rect 11376 16666 11384 16673
rect 11440 16666 11450 16722
rect 11376 16658 11450 16666
rect 10740 16586 10796 16592
rect 10740 16148 10796 16530
rect 10607 15485 10676 15528
rect 10607 5778 10650 15485
rect 10747 15383 10789 16148
rect 29489 15528 29519 17080
rect 29593 17013 29645 17019
rect 29571 16961 29593 17005
rect 29571 16955 29645 16961
rect 29571 15885 29606 16955
rect 29696 16879 29702 16884
rect 29665 16832 29702 16879
rect 29754 16832 29760 16884
rect 29665 16004 29707 16832
rect 29764 16738 29816 16744
rect 29764 16102 29816 16686
rect 29888 16592 29940 16598
rect 29888 16534 29940 16540
rect 29894 16212 29934 16534
rect 29888 16206 29940 16212
rect 29888 16148 29940 16154
rect 29758 16050 29764 16102
rect 29816 16050 29822 16102
rect 29660 15998 29712 16004
rect 29660 15940 29712 15946
rect 29563 15879 29615 15885
rect 29563 15821 29615 15827
rect 30362 15637 30409 34915
rect 30486 28454 30492 28506
rect 30544 28454 30550 28506
rect 30495 15772 30541 28454
rect 30492 15766 30544 15772
rect 30492 15708 30544 15714
rect 30360 15631 30412 15637
rect 30360 15573 30412 15579
rect 29478 15522 29530 15528
rect 29478 15464 29530 15470
rect 10725 15341 10789 15383
rect 10725 5855 10767 15341
rect 13652 15283 13658 15294
rect 10811 15253 13658 15283
rect 10811 5931 10841 15253
rect 13652 15242 13658 15253
rect 13710 15242 13716 15294
rect 13438 15034 14804 15208
rect 17532 15050 17716 15152
rect 17532 14924 17586 15050
rect 17674 14924 17716 15050
rect 17532 14882 17716 14924
rect 11104 13452 11110 13504
rect 11162 13452 11168 13504
rect 11412 13444 11418 13496
rect 11470 13444 11476 13496
rect 11723 13449 11729 13501
rect 11781 13449 11787 13501
rect 12026 13460 12032 13512
rect 12084 13460 12090 13512
rect 12348 13442 12354 13494
rect 12406 13442 12412 13494
rect 12666 13452 12672 13504
rect 12724 13452 12730 13504
rect 12981 13445 12987 13497
rect 13039 13445 13045 13497
rect 13294 13444 13300 13496
rect 13352 13444 13358 13496
rect 17410 11646 17640 11758
rect 17562 11272 17688 11316
rect 17562 11148 17602 11272
rect 17664 11148 17688 11272
rect 17562 11102 17688 11148
rect 10940 9905 11014 10160
rect 10940 9831 12459 9905
rect 12533 9831 13663 9905
rect 12453 9245 12459 9319
rect 12533 9245 12539 9319
rect 11746 7864 11752 7968
rect 11856 7864 11862 7968
rect 13589 7495 13663 9831
rect 29210 8380 29302 8400
rect 29210 8320 29220 8380
rect 29280 8320 29302 8380
rect 29210 8304 29302 8320
rect 13589 7421 13839 7495
rect 13205 6606 13265 6612
rect 13205 6540 13265 6546
rect 10811 5901 12225 5931
rect 10725 5813 12145 5855
rect 10607 5735 12047 5778
rect 12004 3524 12047 5735
rect 12103 3617 12145 5813
rect 12195 4447 12225 5901
rect 12288 5789 12512 5796
rect 12288 5656 12307 5789
rect 12485 5656 12512 5789
rect 12288 5642 12512 5656
rect 12816 4504 12920 4510
rect 12195 4417 12437 4447
rect 12816 4394 12920 4400
rect 13270 4495 13374 4510
rect 13765 4495 13839 7421
rect 17668 7456 17948 7580
rect 17668 7390 17706 7456
rect 17928 7390 17948 7456
rect 17668 7376 17948 7390
rect 13270 4421 13839 4495
rect 13270 4394 13374 4421
rect 14912 3982 15060 4546
rect 20174 4590 20260 4602
rect 20174 4530 20186 4590
rect 20246 4530 20260 4590
rect 20174 4520 20260 4530
rect 23198 4586 23284 4596
rect 23198 4526 23212 4586
rect 23272 4526 23284 4586
rect 23198 4514 23284 4526
rect 26196 4582 26282 4598
rect 26196 4522 26206 4582
rect 26266 4522 26282 4582
rect 26196 4516 26282 4522
rect 23202 3622 23282 3636
rect 23202 3617 23216 3622
rect 12103 3575 23216 3617
rect 23202 3570 23216 3575
rect 23268 3570 23282 3622
rect 23202 3556 23282 3570
rect 29366 3524 29409 4607
rect 12004 3481 29409 3524
<< via1 >>
rect 6686 45044 6746 45050
rect 6686 44996 6692 45044
rect 6692 44996 6740 45044
rect 6740 44996 6746 45044
rect 6686 44990 6746 44996
rect 14970 45030 15022 45082
rect 15520 45008 15572 45060
rect 16066 45016 16118 45068
rect 17726 45036 17778 45088
rect 18258 45022 18344 45098
rect 18834 45012 18886 45064
rect 27616 45014 27668 45066
rect 25176 44806 25236 44866
rect 27336 44811 27388 44863
rect 2706 28758 2826 28878
rect 2712 28078 2832 28198
rect 19198 44396 19252 44448
rect 30078 34878 30198 34998
rect 3132 24704 3214 24780
rect 2738 18538 2790 18590
rect 5590 18538 5642 18590
rect 2598 18410 2650 18462
rect 4302 18410 4354 18462
rect 29524 20804 29576 20856
rect 29514 17080 29566 17132
rect 7520 16526 7576 16582
rect 7520 16222 7576 16278
rect 11384 16666 11440 16722
rect 10740 16530 10796 16586
rect 29593 16961 29645 17013
rect 29702 16832 29754 16884
rect 29764 16686 29816 16738
rect 29888 16540 29940 16592
rect 29888 16154 29940 16206
rect 29764 16050 29816 16102
rect 29660 15946 29712 15998
rect 29563 15827 29615 15879
rect 30492 28454 30544 28506
rect 30492 15714 30544 15766
rect 30360 15579 30412 15631
rect 29478 15470 29530 15522
rect 13658 15242 13710 15294
rect 10972 15066 11060 15162
rect 17586 14924 17674 15050
rect 11110 13452 11162 13504
rect 11418 13444 11470 13496
rect 11729 13449 11781 13501
rect 12032 13460 12084 13512
rect 12354 13442 12406 13494
rect 12672 13452 12724 13504
rect 12987 13445 13039 13497
rect 13300 13444 13352 13496
rect 12324 12534 12588 12680
rect 17232 12143 17293 12204
rect 20204 12130 20264 12190
rect 23182 12134 23242 12194
rect 26216 12126 26276 12186
rect 29196 12120 29292 12218
rect 15710 11610 15964 11720
rect 17602 11148 17664 11272
rect 12459 9831 12533 9905
rect 11010 9542 11256 9654
rect 12459 9245 12533 9319
rect 11752 7864 11856 7968
rect 17214 8346 17274 8406
rect 20192 8338 20252 8398
rect 23220 8330 23280 8390
rect 26224 8342 26284 8402
rect 29220 8320 29280 8380
rect 15678 7818 15938 7920
rect 13205 6546 13265 6606
rect 12314 6006 12600 6126
rect 12307 5656 12485 5789
rect 12816 4400 12920 4504
rect 17706 7390 17928 7456
rect 17188 4540 17248 4600
rect 20186 4530 20246 4590
rect 23212 4526 23272 4586
rect 26206 4522 26266 4582
rect 15670 4018 15930 4120
rect 12312 3676 12640 3804
rect 23216 3570 23268 3622
<< metal2 >>
rect 12734 45092 12828 45112
rect 6660 45050 6774 45076
rect 6660 44990 6686 45050
rect 6746 44990 6774 45050
rect 12734 45032 12750 45092
rect 12810 45032 12828 45092
rect 12734 45008 12828 45032
rect 14382 45062 14476 45130
rect 6660 44962 6774 44990
rect 12766 44862 12794 45008
rect 14382 45002 14404 45062
rect 14464 45002 14476 45062
rect 14382 44976 14476 45002
rect 14928 45086 15070 45118
rect 14928 45026 14966 45086
rect 15026 45026 15070 45086
rect 14928 44988 15070 45026
rect 15490 45064 15606 45094
rect 15490 45004 15516 45064
rect 15576 45004 15606 45064
rect 11458 44834 12794 44862
rect 11458 44674 11486 44834
rect 14407 44779 14461 44976
rect 15490 44972 15606 45004
rect 16038 45072 16146 45100
rect 16038 45012 16062 45072
rect 16122 45012 16146 45072
rect 16038 44976 16146 45012
rect 16594 45062 16700 45088
rect 16594 45002 16618 45062
rect 16678 45002 16700 45062
rect 16594 44976 16700 45002
rect 17128 45066 17280 45114
rect 17128 45006 17162 45066
rect 17222 45006 17280 45066
rect 17704 45092 17808 45124
rect 17704 45032 17722 45092
rect 17782 45032 17808 45092
rect 17704 45012 17808 45032
rect 18244 45098 18370 45124
rect 18244 45022 18258 45098
rect 18344 45022 18370 45098
rect 16627 44811 16668 44976
rect 17128 44956 17280 45006
rect 18244 44988 18370 45022
rect 18796 45068 18910 45088
rect 18796 45008 18830 45068
rect 18890 45008 18910 45068
rect 18796 44982 18910 45008
rect 26490 45080 26668 45106
rect 26490 44988 26516 45080
rect 26608 44988 26668 45080
rect 17164 44825 17219 44956
rect 26490 44942 26668 44988
rect 27062 45088 27204 45116
rect 27062 45028 27098 45088
rect 27158 45028 27204 45088
rect 27062 44982 27204 45028
rect 27596 45070 27686 45084
rect 27596 45010 27612 45070
rect 27672 45010 27686 45070
rect 27596 44994 27686 45010
rect 28186 45066 28286 45088
rect 28186 45006 28206 45066
rect 28266 45006 28286 45066
rect 28186 44984 28286 45006
rect 2398 44646 11486 44674
rect 11613 44725 14461 44779
rect 15006 44770 16668 44811
rect 16768 44784 17219 44825
rect 25160 44866 25256 44880
rect 25160 44806 25176 44866
rect 25236 44806 25256 44866
rect 25160 44796 25256 44806
rect 2398 27694 2426 44646
rect 11613 44571 11667 44725
rect 15006 44664 15047 44770
rect 16780 44735 16821 44784
rect 16852 44770 17219 44784
rect 15106 44702 16821 44735
rect 26516 44734 26608 44942
rect 15106 44694 15860 44702
rect 15980 44694 16821 44702
rect 2493 44517 11667 44571
rect 11743 44623 15054 44664
rect 2493 27937 2547 44517
rect 11743 44472 11784 44623
rect 2915 44431 11784 44472
rect 11865 44581 15054 44582
rect 15106 44581 15147 44694
rect 15890 44664 15950 44673
rect 15890 44595 15950 44604
rect 16908 44642 26608 44734
rect 11865 44540 15147 44581
rect 11865 44529 15054 44540
rect 2700 28878 2840 28884
rect 2700 28758 2706 28878
rect 2826 28758 2840 28878
rect 2700 28750 2840 28758
rect 2630 28198 2844 28214
rect 2630 28078 2712 28198
rect 2832 28078 2844 28198
rect 2630 28070 2844 28078
rect 2493 27883 2801 27937
rect 2398 27666 2646 27694
rect 2459 27202 2519 27211
rect 2459 27133 2519 27142
rect 2469 23885 2508 27133
rect 2618 25870 2646 27666
rect 2747 26113 2801 27883
rect 2915 26283 2978 44431
rect 11865 44380 11918 44529
rect 12760 44462 12854 44478
rect 12760 44402 12774 44462
rect 12834 44402 12854 44462
rect 12760 44382 12854 44402
rect 3070 44327 11918 44380
rect 3070 26442 3123 44327
rect 15906 44302 15934 44595
rect 16908 44354 17000 44642
rect 27100 44532 27156 44982
rect 27310 44867 27430 44882
rect 27310 44807 27332 44867
rect 27392 44807 27430 44867
rect 27310 44786 27430 44807
rect 18978 44482 27156 44532
rect 18978 44476 19164 44482
rect 19290 44476 27156 44482
rect 17932 44384 17988 44432
rect 18978 44384 19034 44476
rect 19192 44448 19258 44454
rect 19192 44396 19198 44448
rect 19252 44396 19258 44448
rect 19192 44390 19258 44396
rect 17932 44328 19034 44384
rect 28222 44370 28250 44984
rect 28222 44342 29514 44370
rect 3194 44064 3203 44124
rect 3263 44117 3272 44124
rect 3263 44070 3381 44117
rect 3263 44064 3272 44070
rect 3334 31915 3381 44070
rect 3297 31868 3381 31915
rect 3297 31680 3344 31868
rect 3184 31612 3372 31680
rect 3070 26389 3400 26442
rect 2915 26220 3028 26283
rect 2747 26059 2863 26113
rect 2618 25842 2710 25870
rect 2682 24102 2710 25842
rect 2809 24303 2863 26059
rect 2965 24545 3028 26220
rect 3096 24780 3236 24796
rect 3096 24704 3132 24780
rect 3214 24704 3236 24780
rect 3096 24676 3236 24704
rect 2965 24482 3092 24545
rect 2809 24249 2959 24303
rect 2682 24074 2778 24102
rect 2459 23442 2517 23885
rect 2420 23433 2556 23442
rect 2420 23323 2433 23433
rect 2543 23323 2556 23433
rect 2420 23312 2556 23323
rect 2750 18596 2778 24074
rect 2905 22098 2959 24249
rect 3029 22413 3092 24482
rect 3029 22350 3290 22413
rect 2905 22078 3150 22098
rect 2872 22073 3150 22078
rect 2872 21963 3013 22073
rect 3123 21963 3150 22073
rect 2872 21958 3150 21963
rect 2940 21944 3150 21958
rect 3219 21409 3290 22350
rect 3045 21402 3293 21409
rect 3003 21398 3293 21402
rect 2998 21393 3293 21398
rect 2998 21283 3003 21393
rect 3113 21339 3293 21393
rect 3113 21303 3289 21339
rect 3113 21283 3198 21303
rect 2998 21278 3198 21283
rect 3003 21274 3113 21278
rect 3347 20738 3400 26389
rect 29486 24928 29514 44342
rect 30078 34998 30198 35004
rect 30078 34872 30198 34878
rect 30244 34313 30386 34326
rect 30244 34203 30261 34313
rect 30371 34203 30386 34313
rect 30244 34188 30386 34203
rect 29746 33633 29882 33638
rect 29746 33523 29756 33633
rect 29866 33523 29882 33633
rect 29746 33508 29882 33523
rect 29790 33049 29832 33508
rect 29707 33007 29832 33049
rect 29560 28846 29662 28860
rect 29560 28790 29582 28846
rect 29638 28790 29662 28846
rect 29560 28770 29662 28790
rect 29486 24900 29564 24928
rect 29536 20862 29564 24900
rect 29595 20954 29626 28770
rect 29595 20923 29657 20954
rect 29524 20856 29576 20862
rect 29524 20798 29576 20804
rect 3322 20516 3424 20738
rect 29502 20692 29580 20708
rect 29502 20636 29512 20692
rect 29568 20636 29580 20692
rect 29502 20612 29580 20636
rect 3322 20468 3434 20516
rect 3324 20462 3434 20468
rect 2738 18590 2790 18596
rect 5584 18538 5590 18590
rect 5642 18538 5648 18590
rect 2738 18532 2790 18538
rect 5602 18512 5630 18538
rect 2582 18466 2666 18478
rect 2582 18406 2594 18466
rect 2654 18406 2666 18466
rect 2582 18394 2666 18406
rect 4294 18462 4362 18470
rect 4294 18410 4302 18462
rect 4354 18410 4362 18462
rect 4294 18404 4362 18410
rect 9450 18426 9510 18435
rect 6890 18218 6918 18368
rect 9450 18357 9510 18366
rect 6965 18218 6974 18234
rect 6890 18190 6974 18218
rect 6965 18174 6974 18190
rect 7034 18174 7043 18234
rect 8784 18110 9002 18124
rect 8784 18050 8806 18110
rect 8866 18050 9002 18110
rect 8784 17996 9002 18050
rect 8146 17938 8284 17954
rect 8146 17878 8162 17938
rect 8222 17878 8284 17938
rect 8146 17864 8284 17878
rect 4942 17788 5002 17797
rect 4942 17719 5002 17728
rect 3001 17384 3010 17444
rect 3070 17384 3079 17444
rect 3636 17170 3728 17182
rect 3636 17110 3654 17170
rect 3714 17110 3728 17170
rect 3636 17098 3728 17110
rect 2368 16256 2424 16622
rect 6232 16398 6288 16654
rect 9452 16646 9508 18357
rect 10072 17616 10324 17636
rect 10072 17556 10094 17616
rect 10154 17556 10324 17616
rect 10072 17536 10324 17556
rect 29525 17138 29555 20612
rect 29514 17132 29566 17138
rect 29514 17074 29566 17080
rect 29626 17013 29657 20923
rect 29587 16961 29593 17013
rect 29645 16971 29657 17013
rect 29645 16961 29651 16971
rect 29707 16890 29749 33007
rect 29832 32953 29968 32962
rect 29832 32843 29845 32953
rect 29955 32843 29968 32953
rect 29832 32832 29968 32843
rect 29702 16884 29754 16890
rect 29702 16826 29754 16832
rect 29874 16738 29926 32832
rect 30293 32439 30339 34188
rect 30293 32393 30541 32439
rect 30218 32273 30354 32284
rect 30218 32163 30233 32273
rect 30343 32246 30354 32273
rect 30343 32190 30440 32246
rect 30343 32163 30354 32190
rect 30218 32154 30354 32163
rect 30247 31593 30347 31602
rect 30024 31508 30247 31568
rect 30024 30434 30084 31508
rect 30247 31474 30347 31483
rect 30138 30913 30274 30924
rect 30138 30803 30153 30913
rect 30263 30803 30274 30913
rect 30138 30794 30274 30803
rect 30034 21156 30074 30434
rect 11376 16722 11450 16732
rect 11376 16666 11384 16722
rect 11440 16666 11450 16722
rect 29758 16686 29764 16738
rect 29816 16686 29926 16738
rect 29966 21116 30074 21156
rect 11376 16658 11450 16666
rect 29966 16620 30006 21116
rect 29932 16592 30006 16620
rect 7520 16582 7576 16588
rect 10734 16530 10740 16586
rect 10796 16530 10802 16586
rect 29882 16540 29888 16592
rect 29940 16546 30006 16592
rect 29940 16540 29946 16546
rect 7520 16520 7576 16526
rect 30190 16474 30226 30794
rect 30384 28370 30440 32190
rect 30495 28512 30541 32393
rect 30492 28506 30544 28512
rect 30492 28448 30544 28454
rect 30384 28314 30478 28370
rect 30301 28193 30357 28202
rect 30301 28074 30357 28083
rect 11118 16438 30226 16474
rect 6232 16342 10836 16398
rect 2368 16200 7358 16256
rect 7514 16222 7520 16278
rect 7576 16222 10704 16278
rect 7302 16160 7358 16200
rect 7302 16104 10558 16160
rect 10502 5694 10558 16104
rect 10648 5816 10704 16222
rect 10780 5926 10836 16342
rect 10944 15162 11076 15184
rect 10944 15066 10972 15162
rect 11060 15066 11076 15162
rect 10944 15042 11076 15066
rect 11118 13510 11154 16438
rect 30311 16400 30347 28074
rect 11426 16364 30347 16400
rect 11110 13504 11162 13510
rect 11426 13502 11462 16364
rect 30422 16314 30478 28314
rect 29662 16309 30478 16314
rect 11732 16264 30478 16309
rect 11732 13507 11777 16264
rect 29662 16258 30478 16264
rect 29882 16200 29888 16206
rect 12038 16160 29888 16200
rect 12038 13518 12078 16160
rect 29882 16154 29888 16160
rect 29940 16154 29946 16206
rect 29764 16102 29816 16108
rect 12354 16050 29764 16102
rect 12032 13512 12084 13518
rect 11110 13446 11162 13452
rect 11418 13496 11470 13502
rect 11418 13438 11470 13444
rect 11729 13501 11781 13507
rect 12032 13454 12084 13460
rect 12354 13494 12406 16050
rect 29764 16044 29816 16050
rect 29654 15993 29660 15998
rect 12677 15951 29660 15993
rect 12677 13510 12719 15951
rect 29654 15946 29660 15951
rect 29712 15946 29718 15998
rect 29557 15871 29563 15879
rect 12995 15836 29563 15871
rect 11729 13443 11781 13449
rect 12672 13504 12724 13510
rect 12995 13503 13030 15836
rect 29557 15827 29563 15836
rect 29615 15827 29621 15879
rect 30486 15763 30492 15766
rect 13303 15717 30492 15763
rect 12672 13446 12724 13452
rect 12987 13497 13039 13503
rect 13303 13502 13349 15717
rect 30486 15714 30492 15717
rect 30544 15714 30550 15766
rect 30354 15629 30360 15631
rect 13549 15582 30360 15629
rect 12354 13436 12406 13442
rect 12987 13439 13039 13445
rect 13300 13496 13352 13502
rect 13300 13438 13352 13444
rect 12296 12680 12626 12708
rect 12296 12534 12324 12680
rect 12588 12534 12626 12680
rect 12296 12506 12626 12534
rect 12459 9905 12533 9911
rect 10968 9654 11296 9688
rect 10968 9542 11010 9654
rect 11256 9542 11296 9654
rect 10968 9504 11296 9542
rect 12459 9319 12533 9831
rect 12459 9239 12533 9245
rect 11752 7968 11856 7974
rect 11752 7664 11856 7864
rect 13196 7769 13205 7829
rect 13265 7822 13274 7829
rect 13549 7822 13596 15582
rect 30354 15579 30360 15582
rect 30412 15579 30418 15631
rect 29472 15511 29478 15522
rect 13669 15481 29478 15511
rect 13669 15300 13699 15481
rect 29472 15470 29478 15481
rect 29530 15470 29536 15522
rect 13658 15294 13710 15300
rect 13658 15236 13710 15242
rect 17562 15050 17688 15066
rect 17562 14924 17586 15050
rect 17674 14924 17688 15050
rect 17562 14898 17688 14924
rect 17186 12204 17338 12260
rect 17186 12143 17232 12204
rect 17293 12143 17338 12204
rect 17186 12114 17338 12143
rect 20158 12190 20310 12230
rect 20158 12130 20204 12190
rect 20264 12130 20310 12190
rect 20158 12084 20310 12130
rect 23142 12194 23294 12238
rect 23142 12134 23182 12194
rect 23242 12134 23294 12194
rect 23142 12092 23294 12134
rect 26160 12186 26312 12236
rect 26160 12126 26216 12186
rect 26276 12126 26312 12186
rect 26160 12090 26312 12126
rect 29162 12218 29324 12230
rect 29162 12120 29196 12218
rect 29292 12120 29324 12218
rect 29162 12100 29324 12120
rect 15688 11720 15994 11742
rect 15688 11610 15710 11720
rect 15964 11610 15994 11720
rect 15688 11592 15994 11610
rect 17562 11272 17688 11316
rect 17562 11148 17602 11272
rect 17664 11148 17688 11272
rect 17562 11102 17688 11148
rect 17158 8406 17310 8444
rect 17158 8346 17214 8406
rect 17274 8346 17310 8406
rect 17158 8298 17310 8346
rect 20162 8398 20314 8456
rect 20162 8338 20192 8398
rect 20252 8338 20314 8398
rect 20162 8310 20314 8338
rect 23172 8390 23324 8456
rect 23172 8330 23220 8390
rect 23280 8330 23324 8390
rect 23172 8310 23324 8330
rect 26176 8402 26328 8454
rect 26176 8342 26224 8402
rect 26284 8342 26328 8402
rect 26176 8308 26328 8342
rect 29210 8380 29302 8400
rect 29210 8320 29220 8380
rect 29280 8320 29302 8380
rect 29210 8304 29302 8320
rect 13265 7775 13596 7822
rect 15648 7920 15954 7944
rect 15648 7818 15678 7920
rect 15938 7818 15954 7920
rect 15648 7794 15954 7818
rect 13265 7769 13274 7775
rect 11752 7560 13860 7664
rect 13199 6604 13205 6606
rect 13265 6604 13271 6606
rect 13198 6548 13205 6604
rect 13265 6548 13272 6604
rect 13199 6546 13205 6548
rect 13265 6546 13271 6548
rect 12290 6126 12620 6152
rect 12290 6006 12314 6126
rect 12600 6006 12620 6126
rect 12290 5984 12620 6006
rect 10780 5870 12200 5926
rect 10648 5760 12050 5816
rect 10502 5638 11908 5694
rect 11852 3364 11908 5638
rect 11994 3472 12050 5760
rect 12144 3588 12200 5870
rect 12288 5789 12512 5796
rect 12288 5656 12307 5789
rect 12485 5656 12512 5789
rect 12288 5642 12512 5656
rect 13756 4504 13860 7560
rect 17674 7456 17940 7466
rect 17674 7390 17706 7456
rect 17928 7390 17940 7456
rect 17674 7376 17940 7390
rect 17174 4600 17260 4612
rect 17174 4540 17188 4600
rect 17248 4540 17260 4600
rect 17174 4530 17260 4540
rect 20174 4590 20260 4602
rect 20174 4530 20186 4590
rect 20246 4530 20260 4590
rect 20174 4520 20260 4530
rect 23198 4586 23284 4596
rect 23198 4526 23212 4586
rect 23272 4526 23284 4586
rect 23198 4514 23284 4526
rect 26196 4582 26282 4598
rect 26196 4522 26206 4582
rect 26266 4522 26282 4582
rect 26196 4516 26282 4522
rect 12810 4400 12816 4504
rect 12920 4400 13860 4504
rect 13756 3950 13860 4400
rect 15646 4120 15962 4142
rect 15646 4018 15670 4120
rect 15930 4018 15962 4120
rect 15646 4002 15962 4018
rect 26795 3950 26958 7765
rect 13756 3945 30517 3950
rect 13710 3792 30517 3945
rect 13767 3787 30517 3792
rect 23202 3626 23282 3636
rect 17179 3588 17188 3590
rect 12144 3532 17188 3588
rect 17179 3530 17188 3532
rect 17248 3530 17257 3590
rect 23202 3566 23212 3626
rect 23272 3566 23282 3626
rect 23202 3556 23282 3566
rect 20177 3472 20186 3474
rect 11994 3416 20186 3472
rect 20177 3414 20186 3416
rect 20246 3414 20255 3474
rect 26197 3364 26206 3366
rect 11852 3308 26206 3364
rect 26197 3306 26206 3308
rect 26266 3306 26275 3366
rect 30354 672 30517 3787
rect 30326 646 30544 672
rect 30326 483 30354 646
rect 30517 483 30544 646
rect 30326 462 30544 483
<< rmetal2 >>
rect 12296 3804 12704 3834
rect 12296 3676 12312 3804
rect 12664 3676 12704 3804
rect 12296 3662 12704 3676
<< via2 >>
rect 6688 44992 6744 45048
rect 12750 45032 12810 45092
rect 14404 45002 14464 45062
rect 14966 45082 15026 45086
rect 14966 45030 14970 45082
rect 14970 45030 15022 45082
rect 15022 45030 15026 45082
rect 14966 45026 15026 45030
rect 15516 45060 15576 45064
rect 15516 45008 15520 45060
rect 15520 45008 15572 45060
rect 15572 45008 15576 45060
rect 15516 45004 15576 45008
rect 16062 45068 16122 45072
rect 16062 45016 16066 45068
rect 16066 45016 16118 45068
rect 16118 45016 16122 45068
rect 16062 45012 16122 45016
rect 16618 45002 16678 45062
rect 17162 45006 17222 45066
rect 17722 45088 17782 45092
rect 17722 45036 17726 45088
rect 17726 45036 17778 45088
rect 17778 45036 17782 45088
rect 17722 45032 17782 45036
rect 18258 45022 18344 45098
rect 18830 45064 18890 45068
rect 18830 45012 18834 45064
rect 18834 45012 18886 45064
rect 18886 45012 18890 45064
rect 18830 45008 18890 45012
rect 26516 44988 26608 45080
rect 27098 45028 27158 45088
rect 27612 45066 27672 45070
rect 27612 45014 27616 45066
rect 27616 45014 27668 45066
rect 27668 45014 27672 45066
rect 27612 45010 27672 45014
rect 28206 45006 28266 45066
rect 25178 44808 25234 44864
rect 15890 44604 15950 44664
rect 2711 28763 2821 28873
rect 2717 28083 2827 28193
rect 2459 27142 2519 27202
rect 12774 44402 12834 44462
rect 27332 44863 27392 44867
rect 27332 44811 27336 44863
rect 27336 44811 27388 44863
rect 27388 44811 27392 44863
rect 27332 44807 27392 44811
rect 3203 44064 3263 44124
rect 3132 24704 3214 24780
rect 2433 23323 2543 23433
rect 3013 21963 3123 22073
rect 3003 21283 3113 21393
rect 30083 34883 30193 34993
rect 30261 34203 30371 34313
rect 29756 33523 29866 33633
rect 29582 28790 29638 28846
rect 29512 20636 29568 20692
rect 2594 18462 2654 18466
rect 2594 18410 2598 18462
rect 2598 18410 2650 18462
rect 2650 18410 2654 18462
rect 2594 18406 2654 18410
rect 9450 18366 9510 18426
rect 6974 18174 7034 18234
rect 8806 18050 8866 18110
rect 8162 17878 8222 17938
rect 4942 17728 5002 17788
rect 3010 17384 3070 17444
rect 3654 17110 3714 17170
rect 10094 17556 10154 17616
rect 29845 32843 29955 32953
rect 30233 32163 30343 32273
rect 30247 31483 30347 31593
rect 30153 30803 30263 30913
rect 30301 28083 30357 28193
rect 10972 15066 11060 15162
rect 12324 12534 12588 12680
rect 11010 9542 11256 9654
rect 13205 7769 13265 7829
rect 17586 14926 17672 15036
rect 17234 12145 17290 12201
rect 20206 12132 20262 12188
rect 23184 12136 23240 12192
rect 26218 12128 26274 12184
rect 29214 12142 29270 12198
rect 15710 11610 15964 11720
rect 17216 8348 17272 8404
rect 20194 8340 20250 8396
rect 23222 8332 23278 8388
rect 26226 8344 26282 8400
rect 29222 8322 29278 8378
rect 15678 7818 15938 7920
rect 13207 6548 13263 6604
rect 12314 6006 12600 6126
rect 12307 5661 12485 5784
rect 17706 7390 17928 7456
rect 17190 4542 17246 4598
rect 20188 4532 20244 4588
rect 23214 4528 23270 4584
rect 26208 4524 26264 4580
rect 15670 4018 15930 4120
rect 12312 3676 12640 3804
rect 12640 3676 12664 3804
rect 17188 3530 17248 3590
rect 23212 3622 23272 3626
rect 23212 3570 23216 3622
rect 23216 3570 23268 3622
rect 23268 3570 23272 3622
rect 23212 3566 23272 3570
rect 20186 3414 20246 3474
rect 26206 3306 26266 3366
rect 30354 483 30517 646
<< metal3 >>
rect 12734 45097 12828 45112
rect 6660 45052 6774 45076
rect 6660 44988 6684 45052
rect 6748 44988 6774 45052
rect 12734 45027 12745 45097
rect 12815 45027 12828 45097
rect 12734 45008 12828 45027
rect 14382 45067 14476 45130
rect 6660 44962 6774 44988
rect 14382 44997 14399 45067
rect 14469 44997 14476 45067
rect 14382 44976 14476 44997
rect 14928 45091 15070 45118
rect 14928 45021 14961 45091
rect 15031 45021 15070 45091
rect 14928 44988 15070 45021
rect 15490 45069 15606 45094
rect 15490 44999 15511 45069
rect 15581 44999 15606 45069
rect 15490 44972 15606 44999
rect 16038 45077 16146 45100
rect 16038 45007 16057 45077
rect 16127 45007 16146 45077
rect 16038 44976 16146 45007
rect 16594 45067 16700 45088
rect 16594 44997 16613 45067
rect 16683 44997 16700 45067
rect 16594 44976 16700 44997
rect 17128 45071 17280 45114
rect 17128 45001 17157 45071
rect 17227 45001 17280 45071
rect 17704 45092 17808 45124
rect 17704 45032 17722 45092
rect 17782 45032 17808 45092
rect 17704 45012 17808 45032
rect 18244 45098 18370 45124
rect 18244 45022 18258 45098
rect 18344 45022 18370 45098
rect 17128 44956 17280 45001
rect 18244 44988 18370 45022
rect 25396 45086 25506 45108
rect 25396 45022 25426 45086
rect 25490 45022 25506 45086
rect 26490 45085 26668 45106
rect 25396 44970 25506 45022
rect 25980 45036 26092 45068
rect 25980 44972 26000 45036
rect 26064 44972 26092 45036
rect 19184 44902 19248 44908
rect 19588 44900 19594 44902
rect 19248 44840 19594 44900
rect 19588 44838 19594 44840
rect 19658 44838 19664 44902
rect 25160 44864 25256 44880
rect 19184 44832 19248 44838
rect 25160 44808 25178 44864
rect 25234 44808 25256 44864
rect 14910 44744 16738 44804
rect 25160 44796 25256 44808
rect 14910 44686 14970 44744
rect 12348 44640 14970 44686
rect 16678 44686 16738 44744
rect 25176 44686 25236 44796
rect 15884 44669 16016 44672
rect 15884 44664 15891 44669
rect 12348 44626 14966 44640
rect 12348 44560 12408 44626
rect 15884 44604 15890 44664
rect 15884 44599 15891 44604
rect 15955 44599 16016 44669
rect 16678 44626 25236 44686
rect 15884 44594 16016 44599
rect 3203 44500 12408 44560
rect 25428 44526 25488 44970
rect 25980 44936 26092 44972
rect 26490 44983 26511 45085
rect 26613 44983 26668 45085
rect 26490 44942 26668 44983
rect 27062 45093 27204 45116
rect 27062 45023 27093 45093
rect 27163 45023 27204 45093
rect 27062 44982 27204 45023
rect 27580 45075 27710 45128
rect 27580 45005 27607 45075
rect 27677 45005 27710 45075
rect 27580 44964 27710 45005
rect 28186 45071 28286 45088
rect 28186 45001 28201 45071
rect 28271 45001 28286 45071
rect 28186 44984 28286 45001
rect 28766 45042 28830 45048
rect 28766 44972 28830 44978
rect 3203 44129 3263 44500
rect 12560 44466 25488 44526
rect 6436 44386 7002 44410
rect 12560 44386 12620 44466
rect 12769 44462 12839 44466
rect 12769 44402 12774 44462
rect 12834 44402 12839 44462
rect 12769 44400 12839 44402
rect 26002 44400 26062 44936
rect 27310 44867 27430 44882
rect 28768 44867 28828 44972
rect 27310 44807 27332 44867
rect 27392 44807 28828 44867
rect 27310 44786 27430 44807
rect 12769 44397 26062 44400
rect 3330 44348 12620 44386
rect 3330 44326 6500 44348
rect 6936 44326 12620 44348
rect 12774 44340 26062 44397
rect 3198 44124 3268 44129
rect 3198 44064 3203 44124
rect 3263 44064 3268 44124
rect 3198 44059 3268 44064
rect 3330 39668 3390 44326
rect 30078 34993 30198 34998
rect 30078 34883 30083 34993
rect 30193 34883 30198 34993
rect 30078 34878 30198 34883
rect 30244 34313 30386 34326
rect 30244 34203 30261 34313
rect 30371 34203 30386 34313
rect 30244 34188 30386 34203
rect 29746 33633 29882 33638
rect 29746 33523 29756 33633
rect 29866 33523 29882 33633
rect 29746 33508 29882 33523
rect 29832 32953 29968 32962
rect 29832 32843 29845 32953
rect 29955 32843 29968 32953
rect 29832 32832 29968 32843
rect 30218 32273 30354 32284
rect 30218 32163 30233 32273
rect 30343 32163 30354 32273
rect 30218 32154 30354 32163
rect 2451 31612 2457 31676
rect 2521 31612 2527 31676
rect 30242 31593 30352 31598
rect 30242 31483 30247 31593
rect 30347 31483 30352 31593
rect 30242 31478 30352 31483
rect 30138 30913 30274 30924
rect 30138 30803 30153 30913
rect 30263 30803 30274 30913
rect 30138 30794 30274 30803
rect 2696 28878 2836 28884
rect 2466 28873 2836 28878
rect 2466 28763 2711 28873
rect 2821 28763 2836 28873
rect 29560 28846 29662 28860
rect 29560 28790 29582 28846
rect 29638 28790 29662 28846
rect 29560 28770 29662 28790
rect 2466 28758 2836 28763
rect 2696 28750 2836 28758
rect 2368 28193 2832 28198
rect 2368 28083 2717 28193
rect 2827 28083 2832 28193
rect 2368 28078 2832 28083
rect 30296 28193 30366 28198
rect 30296 28083 30301 28193
rect 30357 28083 30366 28193
rect 30296 28078 30366 28083
rect 3092 27518 3212 27524
rect 2636 27398 3380 27518
rect 3092 27392 3212 27398
rect 2446 27207 2540 27240
rect 2446 27137 2454 27207
rect 2524 27137 2540 27207
rect 2446 27126 2540 27137
rect 3290 27129 3351 27398
rect 3290 27068 3392 27129
rect 2961 26833 3079 26839
rect 2961 26709 3079 26715
rect 2872 26038 2878 26158
rect 2998 26038 3004 26158
rect 3093 24997 3099 25061
rect 3163 25059 3169 25061
rect 3331 25059 3392 27068
rect 3163 24998 3392 25059
rect 3163 24997 3169 24998
rect 3096 24780 3236 24796
rect 3096 24704 3132 24780
rect 3214 24704 3236 24780
rect 3096 24676 3236 24704
rect 3118 23966 3176 24034
rect 3118 23902 3140 23966
rect 3204 23902 3260 23936
rect 3118 23888 3260 23902
rect 3152 23856 3260 23888
rect 2420 23433 2556 23442
rect 2420 23323 2433 23433
rect 2543 23323 2556 23433
rect 2420 23312 2556 23323
rect 2940 22073 3150 22098
rect 2940 21963 3013 22073
rect 3123 21963 3150 22073
rect 2940 21944 3150 21963
rect 2998 21393 3118 21398
rect 2998 21283 3003 21393
rect 3113 21283 3118 21393
rect 2998 21278 3118 21283
rect 29480 20696 29580 20708
rect 29480 20632 29508 20696
rect 29572 20632 29580 20696
rect 29480 20544 29580 20632
rect 2582 18471 2678 18504
rect 2582 18401 2589 18471
rect 2659 18401 2678 18471
rect 2582 18394 2678 18401
rect 9434 18431 9578 18446
rect 9434 18361 9445 18431
rect 9515 18361 9578 18431
rect 9434 18346 9578 18361
rect 6969 18234 7039 18239
rect 7788 18234 7794 18236
rect 6969 18174 6974 18234
rect 7034 18174 7794 18234
rect 6969 18169 7039 18174
rect 7788 18172 7794 18174
rect 7858 18172 7864 18236
rect 8784 18110 9002 18124
rect 8784 18078 8806 18110
rect 8866 18078 9002 18110
rect 8784 18014 8804 18078
rect 8868 18014 9002 18078
rect 8784 17996 9002 18014
rect 8146 17943 8284 17954
rect 8146 17873 8157 17943
rect 8227 17873 8284 17943
rect 8146 17864 8284 17873
rect 4937 17788 5007 17793
rect 7796 17788 7802 17790
rect 4937 17728 4942 17788
rect 5002 17728 7802 17788
rect 4937 17723 5007 17728
rect 7796 17726 7802 17728
rect 7866 17726 7872 17790
rect 3290 17600 3296 17664
rect 3360 17662 3366 17664
rect 7780 17662 7786 17664
rect 3360 17602 7786 17662
rect 3360 17600 3366 17602
rect 7780 17600 7786 17602
rect 7850 17600 7856 17664
rect 10072 17621 10324 17636
rect 10072 17551 10089 17621
rect 10159 17551 10324 17621
rect 10072 17536 10324 17551
rect 3005 17444 3075 17449
rect 7796 17446 7860 17452
rect 3005 17384 3010 17444
rect 3070 17384 7796 17444
rect 3005 17379 3075 17384
rect 7796 17376 7860 17382
rect 3148 17255 3154 17319
rect 3218 17318 3224 17319
rect 3218 17257 7676 17318
rect 3218 17255 3224 17257
rect 7615 17227 7676 17257
rect 7786 17227 7792 17229
rect 3636 17170 3728 17182
rect 3636 17110 3654 17170
rect 3714 17110 7178 17170
rect 7615 17166 7792 17227
rect 7786 17165 7792 17166
rect 7856 17165 7862 17229
rect 3636 17098 3728 17110
rect 7118 17048 7178 17110
rect 7746 17048 7752 17050
rect 7118 16988 7752 17048
rect 7746 16986 7752 16988
rect 7816 16986 7822 17050
rect 6550 15162 11076 15184
rect 6550 15156 10972 15162
rect 6550 15066 6572 15156
rect 6846 15066 10972 15156
rect 11060 15066 11076 15162
rect 6550 15042 11076 15066
rect 17546 15044 17942 15074
rect 10672 9690 10836 15042
rect 17546 15036 17834 15044
rect 17546 14926 17586 15036
rect 17672 14926 17834 15036
rect 17546 14908 17834 14926
rect 17922 14908 17942 15044
rect 17546 14884 17942 14908
rect 12296 12680 12626 12708
rect 12296 12534 12324 12680
rect 12588 12534 12626 12680
rect 12296 12506 12626 12534
rect 17186 12205 17338 12260
rect 17186 12141 17230 12205
rect 17294 12141 17338 12205
rect 17186 12114 17338 12141
rect 20158 12192 20310 12230
rect 20158 12128 20202 12192
rect 20266 12128 20310 12192
rect 20158 12084 20310 12128
rect 23142 12196 23294 12238
rect 23142 12132 23180 12196
rect 23244 12132 23294 12196
rect 23142 12092 23294 12132
rect 26160 12188 26312 12236
rect 26160 12124 26214 12188
rect 26278 12124 26312 12188
rect 26160 12090 26312 12124
rect 29162 12202 29324 12230
rect 29162 12138 29210 12202
rect 29274 12138 29324 12202
rect 29162 12100 29324 12138
rect 17788 11766 18026 11802
rect 15688 11720 15994 11742
rect 15688 11610 15710 11720
rect 15964 11610 15994 11720
rect 15688 11592 15994 11610
rect 17772 11720 18026 11766
rect 17772 11628 17820 11720
rect 17994 11628 18026 11720
rect 17772 11608 17826 11628
rect 17788 11590 17826 11608
rect 17808 11296 17826 11590
rect 17548 11130 17826 11296
rect 17958 11590 18026 11628
rect 17958 11130 18004 11590
rect 17548 11110 18004 11130
rect 17548 11106 17864 11110
rect 10672 9654 11300 9690
rect 10672 9542 11010 9654
rect 11256 9542 11300 9654
rect 10672 9502 11300 9542
rect 10814 5844 11002 9502
rect 17158 8408 17310 8444
rect 17158 8344 17212 8408
rect 17276 8344 17310 8408
rect 17158 8298 17310 8344
rect 20162 8400 20314 8456
rect 20162 8336 20190 8400
rect 20254 8336 20314 8400
rect 20162 8310 20314 8336
rect 23172 8392 23324 8456
rect 23172 8328 23218 8392
rect 23282 8328 23324 8392
rect 23172 8310 23324 8328
rect 26176 8404 26328 8454
rect 26176 8340 26222 8404
rect 26286 8340 26328 8404
rect 26176 8308 26328 8340
rect 29170 8382 29322 8440
rect 29170 8318 29218 8382
rect 29282 8318 29322 8382
rect 29170 8294 29322 8318
rect 15648 7920 15954 7944
rect 13200 7829 13270 7834
rect 13200 7769 13205 7829
rect 13265 7769 13270 7829
rect 15648 7818 15678 7920
rect 15938 7818 15954 7920
rect 15648 7794 15954 7818
rect 13200 7764 13270 7769
rect 13205 6609 13265 7764
rect 17782 7650 18032 7756
rect 17782 7486 17836 7650
rect 17664 7470 17836 7486
rect 17986 7470 18032 7650
rect 17664 7456 18032 7470
rect 17664 7390 17706 7456
rect 17928 7418 18032 7456
rect 17928 7390 17964 7418
rect 17664 7374 17964 7390
rect 13202 6604 13268 6609
rect 13202 6548 13207 6604
rect 13263 6548 13268 6604
rect 13202 6543 13268 6548
rect 12290 6126 12620 6152
rect 12290 6006 12314 6126
rect 12600 6006 12620 6126
rect 12290 5984 12620 6006
rect 10814 5796 12490 5844
rect 10814 5784 12512 5796
rect 10814 5661 12307 5784
rect 12485 5661 12512 5784
rect 10814 5656 12512 5661
rect 12288 5642 12512 5656
rect 17185 4598 17251 4603
rect 17185 4542 17190 4598
rect 17246 4542 17251 4598
rect 17185 4537 17251 4542
rect 20183 4588 20249 4593
rect 15646 4120 15962 4142
rect 15646 4018 15670 4120
rect 15930 4018 15962 4120
rect 15646 4002 15962 4018
rect 12296 3804 12704 3834
rect 12296 3676 12312 3804
rect 12664 3676 12704 3804
rect 12296 3662 12704 3676
rect 17188 3595 17248 4537
rect 20183 4532 20188 4588
rect 20244 4532 20249 4588
rect 20183 4527 20249 4532
rect 23209 4584 23275 4589
rect 23209 4528 23214 4584
rect 23270 4528 23275 4584
rect 17183 3590 17253 3595
rect 17183 3530 17188 3590
rect 17248 3530 17253 3590
rect 17183 3525 17253 3530
rect 20186 3479 20246 4527
rect 23209 4523 23275 4528
rect 26203 4580 26269 4585
rect 26203 4524 26208 4580
rect 26264 4524 26269 4580
rect 23212 3636 23272 4523
rect 26203 4519 26269 4524
rect 23202 3626 23282 3636
rect 23202 3566 23212 3626
rect 23272 3566 23282 3626
rect 23202 3556 23282 3566
rect 20181 3474 20251 3479
rect 20181 3414 20186 3474
rect 20246 3414 20251 3474
rect 20181 3409 20251 3414
rect 26206 3371 26266 4519
rect 26201 3366 26271 3371
rect 26201 3306 26206 3366
rect 26266 3306 26271 3366
rect 26201 3301 26271 3306
rect 30326 651 30544 672
rect 30326 478 30349 651
rect 30522 478 30544 651
rect 30326 462 30544 478
<< rmetal3 >>
rect 18796 45068 18910 45088
rect 18796 45008 18830 45068
rect 18890 45008 18910 45068
rect 18796 44982 18910 45008
<< via3 >>
rect 6684 45048 6748 45052
rect 6684 44992 6688 45048
rect 6688 44992 6744 45048
rect 6744 44992 6748 45048
rect 6684 44988 6748 44992
rect 12745 45092 12815 45097
rect 12745 45032 12750 45092
rect 12750 45032 12810 45092
rect 12810 45032 12815 45092
rect 12745 45027 12815 45032
rect 14399 45062 14469 45067
rect 14399 45002 14404 45062
rect 14404 45002 14464 45062
rect 14464 45002 14469 45062
rect 14399 44997 14469 45002
rect 14961 45086 15031 45091
rect 14961 45026 14966 45086
rect 14966 45026 15026 45086
rect 15026 45026 15031 45086
rect 14961 45021 15031 45026
rect 15511 45064 15581 45069
rect 15511 45004 15516 45064
rect 15516 45004 15576 45064
rect 15576 45004 15581 45064
rect 15511 44999 15581 45004
rect 16057 45072 16127 45077
rect 16057 45012 16062 45072
rect 16062 45012 16122 45072
rect 16122 45012 16127 45072
rect 16057 45007 16127 45012
rect 16613 45062 16683 45067
rect 16613 45002 16618 45062
rect 16618 45002 16678 45062
rect 16678 45002 16683 45062
rect 16613 44997 16683 45002
rect 17157 45066 17227 45071
rect 17157 45006 17162 45066
rect 17162 45006 17222 45066
rect 17222 45006 17227 45066
rect 17157 45001 17227 45006
rect 25426 45022 25490 45086
rect 26000 44972 26064 45036
rect 19184 44838 19248 44902
rect 19594 44838 19658 44902
rect 15891 44664 15955 44669
rect 15891 44604 15950 44664
rect 15950 44604 15955 44664
rect 15891 44599 15955 44604
rect 26511 45080 26613 45085
rect 26511 44988 26516 45080
rect 26516 44988 26608 45080
rect 26608 44988 26613 45080
rect 26511 44983 26613 44988
rect 27093 45088 27163 45093
rect 27093 45028 27098 45088
rect 27098 45028 27158 45088
rect 27158 45028 27163 45088
rect 27093 45023 27163 45028
rect 27607 45070 27677 45075
rect 27607 45010 27612 45070
rect 27612 45010 27672 45070
rect 27672 45010 27677 45070
rect 27607 45005 27677 45010
rect 28201 45066 28271 45071
rect 28201 45006 28206 45066
rect 28206 45006 28266 45066
rect 28266 45006 28271 45066
rect 28201 45001 28271 45006
rect 28766 44978 28830 45042
rect 2457 31612 2521 31676
rect 2454 27202 2524 27207
rect 2454 27142 2459 27202
rect 2459 27142 2519 27202
rect 2519 27142 2524 27202
rect 2454 27137 2524 27142
rect 2961 26715 3079 26833
rect 2878 26038 2998 26158
rect 3099 24997 3163 25061
rect 3140 23902 3204 23966
rect 29508 20692 29572 20696
rect 29508 20636 29512 20692
rect 29512 20636 29568 20692
rect 29568 20636 29572 20692
rect 29508 20632 29572 20636
rect 2589 18466 2659 18471
rect 2589 18406 2594 18466
rect 2594 18406 2654 18466
rect 2654 18406 2659 18466
rect 2589 18401 2659 18406
rect 9445 18426 9515 18431
rect 9445 18366 9450 18426
rect 9450 18366 9510 18426
rect 9510 18366 9515 18426
rect 9445 18361 9515 18366
rect 7794 18172 7858 18236
rect 8804 18050 8806 18078
rect 8806 18050 8866 18078
rect 8866 18050 8868 18078
rect 8804 18014 8868 18050
rect 8157 17938 8227 17943
rect 8157 17878 8162 17938
rect 8162 17878 8222 17938
rect 8222 17878 8227 17938
rect 8157 17873 8227 17878
rect 7802 17726 7866 17790
rect 3296 17600 3360 17664
rect 7786 17600 7850 17664
rect 10089 17616 10159 17621
rect 10089 17556 10094 17616
rect 10094 17556 10154 17616
rect 10154 17556 10159 17616
rect 10089 17551 10159 17556
rect 7796 17382 7860 17446
rect 3154 17255 3218 17319
rect 7792 17165 7856 17229
rect 7752 16986 7816 17050
rect 6572 15066 6846 15156
rect 17834 14908 17922 15044
rect 12324 12534 12588 12680
rect 17230 12201 17294 12205
rect 17230 12145 17234 12201
rect 17234 12145 17290 12201
rect 17290 12145 17294 12201
rect 17230 12141 17294 12145
rect 20202 12188 20266 12192
rect 20202 12132 20206 12188
rect 20206 12132 20262 12188
rect 20262 12132 20266 12188
rect 20202 12128 20266 12132
rect 23180 12192 23244 12196
rect 23180 12136 23184 12192
rect 23184 12136 23240 12192
rect 23240 12136 23244 12192
rect 23180 12132 23244 12136
rect 26214 12184 26278 12188
rect 26214 12128 26218 12184
rect 26218 12128 26274 12184
rect 26274 12128 26278 12184
rect 26214 12124 26278 12128
rect 29210 12198 29274 12202
rect 29210 12142 29214 12198
rect 29214 12142 29270 12198
rect 29270 12142 29274 12198
rect 29210 12138 29274 12142
rect 15710 11610 15964 11720
rect 17820 11628 17994 11720
rect 17826 11130 17958 11628
rect 17212 8404 17276 8408
rect 17212 8348 17216 8404
rect 17216 8348 17272 8404
rect 17272 8348 17276 8404
rect 17212 8344 17276 8348
rect 20190 8396 20254 8400
rect 20190 8340 20194 8396
rect 20194 8340 20250 8396
rect 20250 8340 20254 8396
rect 20190 8336 20254 8340
rect 23218 8388 23282 8392
rect 23218 8332 23222 8388
rect 23222 8332 23278 8388
rect 23278 8332 23282 8388
rect 23218 8328 23282 8332
rect 26222 8400 26286 8404
rect 26222 8344 26226 8400
rect 26226 8344 26282 8400
rect 26282 8344 26286 8400
rect 26222 8340 26286 8344
rect 29218 8378 29282 8382
rect 29218 8322 29222 8378
rect 29222 8322 29278 8378
rect 29278 8322 29282 8378
rect 29218 8318 29282 8322
rect 15678 7818 15938 7920
rect 17836 7470 17986 7650
rect 12314 6006 12600 6126
rect 15670 4018 15930 4120
rect 12312 3676 12664 3804
rect 30349 646 30522 651
rect 30349 483 30354 646
rect 30354 483 30517 646
rect 30517 483 30522 646
rect 30349 478 30522 483
<< metal4 >>
rect 6134 45040 6194 45152
rect 6686 45076 6746 45152
rect 6660 45052 6774 45076
rect 6660 45040 6684 45052
rect 6134 44988 6684 45040
rect 6748 45040 6774 45052
rect 7238 45040 7298 45152
rect 7790 45040 7850 45152
rect 8342 45040 8402 45152
rect 8894 45040 8954 45152
rect 9446 45040 9506 45152
rect 9998 45040 10058 45152
rect 10550 45040 10610 45152
rect 11102 45040 11162 45152
rect 11654 45040 11714 45152
rect 6748 44988 11714 45040
rect 6134 44980 11714 44988
rect 6134 44952 6194 44980
rect 6660 44962 6774 44980
rect 6686 44952 6746 44962
rect 7238 44952 7298 44980
rect 7790 44952 7850 44980
rect 8342 44952 8402 44980
rect 8894 44952 8954 44980
rect 9446 44952 9506 44980
rect 9998 44952 10058 44980
rect 10550 44952 10610 44980
rect 11102 44952 11162 44980
rect 11654 44952 11714 44980
rect 12206 45038 12266 45152
rect 12758 45112 12818 45152
rect 12734 45097 12828 45112
rect 12206 44952 12274 45038
rect 12734 45027 12745 45097
rect 12815 45027 12828 45097
rect 13310 45089 13370 45152
rect 12734 45008 12828 45027
rect 12758 44952 12818 45008
rect 13304 44952 13370 45089
rect 13862 45068 13922 45152
rect 14414 45130 14474 45152
rect 12214 44862 12274 44952
rect 2594 44802 12274 44862
rect 2456 31676 2522 31677
rect 2456 31612 2457 31676
rect 2521 31612 2522 31676
rect 2456 31611 2522 31612
rect 2459 27228 2519 31611
rect 2446 27207 2532 27228
rect 2446 27137 2454 27207
rect 2524 27137 2532 27207
rect 2446 27126 2532 27137
rect 2594 18478 2654 44802
rect 13304 44707 13367 44952
rect 3412 44682 13367 44707
rect 2948 44644 13367 44682
rect 2948 44612 3475 44644
rect 2948 44608 3012 44612
rect 2948 26985 3011 44608
rect 13824 44552 13944 45068
rect 14382 45067 14476 45130
rect 14966 45118 15026 45152
rect 14382 44997 14399 45067
rect 14469 44997 14476 45067
rect 14382 44976 14476 44997
rect 14928 45091 15070 45118
rect 15518 45094 15578 45152
rect 16070 45100 16130 45152
rect 14928 45021 14961 45091
rect 15031 45021 15070 45091
rect 14928 44988 15070 45021
rect 15490 45069 15606 45094
rect 15490 44999 15511 45069
rect 15581 44999 15606 45069
rect 14414 44952 14474 44976
rect 14966 44952 15026 44988
rect 15490 44972 15606 44999
rect 16038 45077 16146 45100
rect 16622 45088 16682 45152
rect 17174 45108 17234 45152
rect 17726 45124 17786 45152
rect 18278 45124 18338 45152
rect 16038 45007 16057 45077
rect 16127 45007 16146 45077
rect 16038 44976 16146 45007
rect 16594 45067 16700 45088
rect 16594 44997 16613 45067
rect 16683 44997 16700 45067
rect 16594 44976 16700 44997
rect 17128 45071 17280 45108
rect 17128 45001 17157 45071
rect 17227 45001 17280 45071
rect 17704 45012 17808 45124
rect 15518 44952 15578 44972
rect 16070 44952 16130 44976
rect 16622 44952 16682 44976
rect 17128 44950 17280 45001
rect 17726 44952 17786 45012
rect 18244 44988 18370 45124
rect 18830 45088 18890 45152
rect 19382 45112 19442 45152
rect 19934 45112 19994 45152
rect 20486 45112 20546 45152
rect 21038 45112 21098 45152
rect 21590 45112 21650 45152
rect 22142 45112 22202 45152
rect 22694 45112 22754 45152
rect 23246 45112 23306 45152
rect 18278 44952 18338 44988
rect 18796 44982 18910 45088
rect 19380 45052 23306 45112
rect 18830 44952 18890 44982
rect 19380 44952 19442 45052
rect 19934 44952 19994 45052
rect 20486 44952 20546 45052
rect 21038 44952 21098 45052
rect 21590 44952 21650 45052
rect 22142 44952 22202 45052
rect 22694 44952 22754 45052
rect 23246 44952 23306 45052
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 45108 25514 45152
rect 25396 45086 25514 45108
rect 25396 45022 25426 45086
rect 25490 45022 25514 45086
rect 26006 45068 26066 45152
rect 26558 45106 26618 45152
rect 27110 45116 27170 45152
rect 26490 45085 26668 45106
rect 25396 44970 25514 45022
rect 25454 44952 25514 44970
rect 25980 45036 26092 45068
rect 25980 44972 26000 45036
rect 26064 44972 26092 45036
rect 19183 44902 19249 44903
rect 19183 44838 19184 44902
rect 19248 44838 19249 44902
rect 19183 44837 19249 44838
rect 15884 44669 15956 44672
rect 15884 44600 15891 44669
rect 15890 44599 15891 44600
rect 15955 44664 15956 44669
rect 19186 44664 19246 44837
rect 15955 44604 19246 44664
rect 15955 44599 15956 44604
rect 15890 44598 15956 44599
rect 2767 26980 3011 26985
rect 2766 26922 3011 26980
rect 3092 44432 13944 44552
rect 2766 26223 2835 26922
rect 3092 26834 3212 44432
rect 6558 42260 6880 44304
rect 2960 26833 3212 26834
rect 2960 26715 2961 26833
rect 3079 26715 3212 26833
rect 2960 26714 3212 26715
rect 2766 26181 2903 26223
rect 2759 26159 2903 26181
rect 2759 26158 2999 26159
rect 2759 26115 2878 26158
rect 2763 26059 2878 26115
rect 2877 26038 2878 26059
rect 2998 26038 2999 26158
rect 2877 26037 2999 26038
rect 3098 25061 3164 25062
rect 3098 25060 3099 25061
rect 2952 24999 3099 25060
rect 2952 23793 3013 24999
rect 3098 24997 3099 24999
rect 3163 24997 3164 25061
rect 3098 24996 3164 24997
rect 3139 23966 3205 23967
rect 3139 23902 3140 23966
rect 3204 23964 3205 23966
rect 3204 23904 3358 23964
rect 3204 23902 3205 23904
rect 3139 23901 3205 23902
rect 2952 23732 3216 23793
rect 2582 18471 2666 18478
rect 2582 18401 2589 18471
rect 2659 18401 2666 18471
rect 2582 18394 2666 18401
rect 3155 17320 3216 23732
rect 3298 17665 3358 23904
rect 3295 17664 3361 17665
rect 3295 17600 3296 17664
rect 3360 17600 3361 17664
rect 3295 17599 3361 17600
rect 3153 17319 3219 17320
rect 3153 17255 3154 17319
rect 3218 17255 3219 17319
rect 3153 17254 3219 17255
rect 6552 15156 6880 42260
rect 7218 44138 7536 44302
rect 19380 44138 19440 44952
rect 25980 44936 26092 44972
rect 26490 44983 26511 45085
rect 26613 44983 26668 45085
rect 26490 44942 26668 44983
rect 27062 45093 27204 45116
rect 27062 45023 27093 45093
rect 27163 45023 27204 45093
rect 27062 44982 27204 45023
rect 27574 45075 27722 45152
rect 28214 45088 28274 45152
rect 27574 45005 27607 45075
rect 27677 45005 27722 45075
rect 27110 44952 27170 44982
rect 27574 44952 27722 45005
rect 28186 45071 28286 45088
rect 28186 45001 28201 45071
rect 28271 45001 28286 45071
rect 28766 45043 28826 45152
rect 28186 44984 28286 45001
rect 28765 45042 28831 45043
rect 28214 44952 28274 44984
rect 28765 44978 28766 45042
rect 28830 44978 28831 45042
rect 28765 44977 28831 44978
rect 28766 44952 28826 44977
rect 29318 44952 29378 45152
rect 19593 44902 19659 44903
rect 19593 44838 19594 44902
rect 19658 44838 19659 44902
rect 19593 44837 19659 44838
rect 19596 44424 19656 44837
rect 19596 44364 29538 44424
rect 7218 44078 19440 44138
rect 7218 15588 7536 44078
rect 29478 20708 29538 44364
rect 29478 20696 29580 20708
rect 29478 20634 29508 20696
rect 29502 20632 29508 20634
rect 29572 20632 29580 20696
rect 29502 20612 29580 20632
rect 9444 18431 9516 18432
rect 9444 18361 9445 18431
rect 9515 18426 9516 18431
rect 9515 18366 29536 18426
rect 9515 18361 9516 18366
rect 9444 18360 9516 18361
rect 7793 18236 7859 18237
rect 7793 18172 7794 18236
rect 7858 18234 7859 18236
rect 7858 18174 28924 18234
rect 7858 18172 7859 18174
rect 7793 18171 7859 18172
rect 8784 18078 9002 18114
rect 8784 18014 8804 18078
rect 8868 18076 9002 18078
rect 8868 18016 26276 18076
rect 8868 18014 9002 18016
rect 8784 18002 9002 18014
rect 8156 17943 8228 17944
rect 8156 17873 8157 17943
rect 8227 17938 8228 17943
rect 8227 17878 25728 17938
rect 8227 17873 8228 17878
rect 8156 17872 8228 17873
rect 7801 17790 7867 17791
rect 7801 17726 7802 17790
rect 7866 17788 7867 17790
rect 7866 17728 23242 17788
rect 7866 17726 7867 17728
rect 7801 17725 7867 17726
rect 7785 17664 7851 17665
rect 7785 17600 7786 17664
rect 7850 17662 7851 17664
rect 7850 17602 9754 17662
rect 7850 17600 7851 17602
rect 7785 17599 7851 17600
rect 9694 17468 9754 17602
rect 10088 17621 10160 17622
rect 10088 17551 10089 17621
rect 10159 17616 10160 17621
rect 10159 17556 22774 17616
rect 10159 17551 10160 17556
rect 10088 17550 10160 17551
rect 7795 17446 7861 17447
rect 7795 17382 7796 17446
rect 7860 17444 7861 17446
rect 7860 17384 9480 17444
rect 9694 17408 20264 17468
rect 7860 17382 7861 17384
rect 7795 17381 7861 17382
rect 9420 17322 9480 17384
rect 9420 17262 19964 17322
rect 7791 17229 7857 17230
rect 7791 17165 7792 17229
rect 7856 17228 7857 17229
rect 7856 17183 9346 17228
rect 7856 17167 17292 17183
rect 7856 17165 7857 17167
rect 7791 17164 7857 17165
rect 9285 17122 17292 17167
rect 7751 17050 7817 17051
rect 7751 16986 7752 17050
rect 7816 17048 7817 17050
rect 7816 16988 16790 17048
rect 7816 16986 7817 16988
rect 7751 16985 7817 16986
rect 7216 15548 7536 15588
rect 6552 15066 6572 15156
rect 6846 15066 6880 15156
rect 6552 2318 6880 15066
rect 7214 4049 7536 15548
rect 12293 12680 12615 12729
rect 12293 12534 12324 12680
rect 12588 12534 12615 12680
rect 12293 6126 12615 12534
rect 15688 11729 15994 11742
rect 12293 6006 12314 6126
rect 12600 6006 12615 6126
rect 12293 4049 12615 6006
rect 15641 11720 15994 11729
rect 15641 11610 15710 11720
rect 15964 11610 15994 11720
rect 15641 11592 15994 11610
rect 15641 7920 15963 11592
rect 16730 8406 16790 16988
rect 17231 12260 17292 17122
rect 17784 15044 18032 15302
rect 17784 14908 17834 15044
rect 17922 14908 18032 15044
rect 17186 12205 17338 12260
rect 17186 12141 17230 12205
rect 17294 12141 17338 12205
rect 17186 12114 17338 12141
rect 17784 11720 18032 14908
rect 17784 11628 17820 11720
rect 17994 11628 18032 11720
rect 17784 11130 17826 11628
rect 17958 11130 18032 11628
rect 17158 8408 17310 8444
rect 17158 8406 17212 8408
rect 16730 8346 17212 8406
rect 17158 8344 17212 8346
rect 17276 8344 17310 8408
rect 17158 8298 17310 8344
rect 15641 7818 15678 7920
rect 15938 7818 15963 7920
rect 15641 4120 15963 7818
rect 17784 7756 18032 11130
rect 19904 8398 19964 17262
rect 20204 12230 20264 17408
rect 20158 12192 20310 12230
rect 20158 12128 20202 12192
rect 20266 12128 20310 12192
rect 20158 12084 20310 12128
rect 20162 8400 20314 8456
rect 20162 8398 20190 8400
rect 19904 8338 20190 8398
rect 20162 8336 20190 8338
rect 20254 8336 20314 8400
rect 20162 8310 20314 8336
rect 22714 8390 22774 17556
rect 23182 12197 23242 17728
rect 23179 12196 23245 12197
rect 23179 12132 23180 12196
rect 23244 12132 23245 12196
rect 23179 12131 23245 12132
rect 23172 8392 23324 8456
rect 23172 8390 23218 8392
rect 22714 8330 23218 8390
rect 23172 8328 23218 8330
rect 23282 8328 23324 8392
rect 25668 8402 25728 17878
rect 26216 12189 26276 18016
rect 26213 12188 26279 12189
rect 26213 12124 26214 12188
rect 26278 12124 26279 12188
rect 26213 12123 26279 12124
rect 26176 8404 26328 8454
rect 26176 8402 26222 8404
rect 25668 8342 26222 8402
rect 23172 8310 23324 8328
rect 26176 8340 26222 8342
rect 26286 8340 26328 8404
rect 26176 8308 26328 8340
rect 28864 8380 28924 18174
rect 29162 12202 29324 12230
rect 29162 12138 29210 12202
rect 29274 12200 29324 12202
rect 29476 12200 29536 18366
rect 29274 12140 29536 12200
rect 29274 12138 29324 12140
rect 29162 12100 29324 12138
rect 29210 8382 29302 8400
rect 29210 8380 29218 8382
rect 28864 8320 29218 8380
rect 29210 8318 29218 8320
rect 29282 8318 29302 8382
rect 29210 8304 29302 8318
rect 17782 7650 18032 7756
rect 17782 7470 17836 7650
rect 17986 7470 18032 7650
rect 17782 7418 18032 7470
rect 15641 4049 15670 4120
rect 7214 4018 15670 4049
rect 15930 4049 15963 4120
rect 15930 4018 16649 4049
rect 7214 3804 16649 4018
rect 7214 3727 12312 3804
rect 6552 1654 6874 2318
rect 6552 1410 6878 1654
rect 7214 1410 7536 3727
rect 12296 3676 12312 3727
rect 12664 3727 16649 3804
rect 12664 3676 12704 3727
rect 12296 3662 12704 3676
rect 6512 1010 6912 1410
rect 7184 1010 7584 1410
rect 6552 720 6878 1010
rect 6552 274 6874 720
rect 7214 314 7536 1010
rect 30326 651 30544 672
rect 30326 478 30349 651
rect 30522 478 30544 651
rect 30326 462 30544 478
rect 7214 274 7534 314
rect 30354 200 30517 462
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 0 26678 200
rect 30354 45 30542 200
rect 30362 0 30542 45
use compr  compr_0
timestamp 1730635755
transform 1 0 9678 0 1 6382
box 1230 -398 4034 3312
use flash_adc2  flash_adc2_0
timestamp 1730635755
transform 1 0 27580 0 1 3786
box -13594 198 2206 11530
use main  main_0
timestamp 1730493024
transform 1 0 2350 0 1 16510
box -4 0 28201 27950
use pass_gate2  pass_gate2_0
timestamp 1730493024
transform 1 0 10882 0 1 4780
box 1380 -1118 2522 1056
use r2r_dac  r2r_dac_0
timestamp 1730635755
transform 1 0 9898 0 1 15400
box 1000 -5458 3772 -192
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 1 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 2 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 3 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 4 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 5 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 6 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 7 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 8 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 9 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 11 nsew signal input
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 12 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 13 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 14 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 15 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 16 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 17 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 18 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 19 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 20 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 21 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 22 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 23 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 24 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 25 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 26 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 27 nsew signal output
flabel metal4 s 6512 1010 6912 1410 0 FreeSans 480 90 0 0 VDPWR
port 28 nsew signal output
flabel metal4 s 7184 1010 7584 1410 0 FreeSans 480 90 0 0 VGND
port 10 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
